module tb;
reg signed [3:0]a;
initial begin
a= 4'b1001;
$display(a);
end
endmodule
