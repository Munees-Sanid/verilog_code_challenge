module tast_name(

)


integer i;
module
task
