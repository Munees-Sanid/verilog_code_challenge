module serial(
	input a,b,
	output y);
assign
