module (
input a,b,c,
output f)
always@(posedge clk)
