module tast_name(

)

task
