module tb;
signed reg[7:0]a;
initial begin
a=-7;
$display("a = %0d",a);
end
endmodule
