module tast_name(

)


integer i;
task
