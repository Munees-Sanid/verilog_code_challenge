module demux(
input a, 
output c,d,e);
