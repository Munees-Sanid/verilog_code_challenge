// simple real time clock 

module rtc(
	input 
