// design code for fsm 

module fsm(
	input
